// slon01.v
module slon01;
endmodule 
//------------------------------------------------------------------------------
//  project:       slon5_test
//  module:        slon5_test
//
//  description:   slon5 start-up
//------------------------------------------------------------------------------

`include "slon5.svh"    

//******************************************************************************
//******************************************************************************
module slon5_test import slon5_pkg::*;
(
    input  logic  ref_clk,
                                 
    input  Dnum_t sw,

    output Dout_t dout,
    output Dnum_t dnum
);

//==============================================================================
//    Settings
//==============================================================================

//==============================================================================
//    Types
//==============================================================================

//==============================================================================
//    Objects
//==============================================================================

logic clk;
logic rst;

//==============================================================================
//     Logic
//==============================================================================

//==============================================================================
//    Instances
//==============================================================================

//------------------------------------------------------------------------------
//    Reset
//------------------------------------------------------------------------------
rst_m rst_inst
(
    .clk ( clk ),
    .q   ( rst )
);

//------------------------------------------------------------------------------
//    pll
//------------------------------------------------------------------------------
`ifndef SIMULATOR
    //---- PLL instance
    pll pll_inst
    (
        .clk_in1  ( ref_clk ),
        .clk_out1 ( clk     )
    );
`else
    assign clk = ref_clk;
`endif


//------------------------------------------------------------------------------
//    slon5_m
//------------------------------------------------------------------------------

slon5_m slon5
(
    .clk  ( clk     ),
    .rst  ( rst     ),
    
    .sw   ( sw      ),
    
    .dout ( dout    ),
    .dnum ( dnum    )
);

//==============================================================================
//    snippets
//==============================================================================

//------------------------------------------------------------------------------
//    SIMULATOR

`ifndef SIMULATOR
    // ***
`else
    // ***
`endif

endmodule : slon5_test


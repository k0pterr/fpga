// slon11.v
module slon11;
endmodule

//------------------------------------------------------------------------------
//  project:       slon5_test
//  module:        slon5_test
//
//  description:   slon5 start-up
//------------------------------------------------------------------------------

`include "slon5.svh"    

//******************************************************************************
//******************************************************************************
module slon5_test import slon5_pkg::*;
(
    input  logic  ref_clk,
                                 
    input  Dnum_t sw,

    output Dout_t dout,
    output Dnum_t dnum
);

//==============================================================================
//    Settings
//==============================================================================

//==============================================================================
//    Types
//==============================================================================

//==============================================================================
//    Objects
//==============================================================================

//==============================================================================
//     Logic
//==============================================================================

//==============================================================================
//    Instances
//==============================================================================

//------------------------------------------------------------------------------
//    slon5_m
//------------------------------------------------------------------------------

slon5_m slon5
(
    .clk  ( 1'bx    ),
    
    .sw   ( sw      ),
    
    .dout ( dout    ),
    .dnum ( dnum    )
);

//==============================================================================
//    snippets
//==============================================================================

//------------------------------------------------------------------------------
//    SIMULATOR

`ifndef SIMULATOR
    // ***
`else
    // ***
`endif

endmodule : slon5_test


//-------------------------------------------------------------------------------
//
//     Project: Any
//
//     Purpose: Default top-level file
//
//
//-------------------------------------------------------------------------------

module top
(
    input  in;
    output out;
);

assign out = in;

endmodule
//-------------------------------------------------------------------------------

// slon21.v
module slon21;
endmodule
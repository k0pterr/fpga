// slon12.sv
module slon12;
endmodule

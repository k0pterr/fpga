//------------------------------------------------------------------------------
//  project:       slon5_test
//  module:        slon5_test
//
//  description:   slon5 start-up
//------------------------------------------------------------------------------

`include "slon5.svh"    

//******************************************************************************
//******************************************************************************
module slon5_test import slon5_pkg::*;
(
`ifdef DIFF_REFCLK
    input  logic  ref_clk_p,
    input  logic  ref_clk_n,
`else
    input  logic  ref_clk,
`endif
                                 
    input  Dnum_t sw,

    output Dout_t dout,
    output Dnum_t dnum
);

//==============================================================================
//    Settings
//==============================================================================

//==============================================================================
//    Types
//==============================================================================

//==============================================================================
//    Objects
//==============================================================================

`ifdef DIFF_REFCLK
logic ref_clk;
`endif

logic clk;
logic rst;

logic pll_locked;

//==============================================================================
//     Logic
//==============================================================================

//==============================================================================
//    Instances
//==============================================================================

//------------------------------------------------------------------------------
//    Reset
//------------------------------------------------------------------------------
rst_m rst_inst
(
    .clk ( clk ),
    .q   ( rst )
);

//------------------------------------------------------------------------------
//    Clock
//------------------------------------------------------------------------------
`ifdef DIFF_REFCLK
IBUFDS diff_clk_200 
(
    .I  ( ref_clk_p ),
    .IB ( ref_clk_n ),
    .O  ( ref_clk   )
);
`endif

pll pll_inst
(
    .clk_in1  ( ref_clk    ),
    .clk_out1 ( clk        ),
    .locked   ( pll_locked )
);
`ifndef SIMULATOR
    //---- PLL instance
`else
//    assign clk = ref_clk;
`endif


//------------------------------------------------------------------------------
//    slon5_m
//------------------------------------------------------------------------------

slon5_m slon5
(
    .clk  ( clk     ),
    .rst  ( rst     ),
    
    .sw   ( sw      ),
    
    .dout ( dout    ),
    .dnum ( dnum    )
);

//==============================================================================
//    snippets
//==============================================================================

//------------------------------------------------------------------------------
//    SIMULATOR

`ifndef SIMULATOR
    // ***
`else
    // ***
`endif

endmodule : slon5_test


//------------------------------------------------------------------------------
//  project:       slon5_test
//  module:        slon5_tb
//
//  description:   slon5 start-up
//------------------------------------------------------------------------------

`include "common.pkg"
`include "slon5.svh"    
`include "slon5_debug.svh"    

           
//******************************************************************************
//******************************************************************************
module slon5_tb import slon5_pkg::*,
                       slon5_generated_pkg::*,
                       slon5_debug_pkg::*;
();

//==============================================================================
//    Settings
//==============================================================================
                               
//------------------------------------------------------------------------------
`define CLK_HALF_PERIOD     5ns
`define WATCH_DOG_TIME   1000ns

//------------------------------------------------------------------------------
parameter real SCALE_MHz = 1e6;
parameter real SCALE_uS  = 1e-6;
parameter real SCALE_nS  = 1e-9;

parameter int SYSTEM_CLOCK  = ((1.0/(`CLK_HALF_PERIOD*2.0*SCALE_nS))/SCALE_MHz);

//==============================================================================
//    Types
//==============================================================================

//==============================================================================
//    Objects
//==============================================================================

bit   clk;
bit   rst;

string sInfo = "slon5_test";

var Dnum_t sw;
var Dnum_t dnum;
var Dout_t dout;

//==============================================================================
//     Logic
//==============================================================================


//------------------------------------------------------------------------------
initial begin  : input_clk
    fork
        begin
            wait (clk == 1);
            wait (clk == 0);
            #200ps;
            rst = 0;
        end
        begin
            rst = 1;
            clk = 0;
            #3000ps;
            forever #`CLK_HALF_PERIOD clk = ~clk;
        end
    join  
end : input_clk

//------------------------------------------------------------------------------
initial begin : stop_WatchDog
    $write("----------------------------------------------------------------\n");
    $write("Simulation start\n");
    $write("----------------------------------------------------------------\n");
    #`WATCH_DOG_TIME
    sInfo = "slon5_test_stop";
    #50ns
    $write("----------------------------------------------------------------\n");
    $write("Simulation stop\n");
    $write("----------------------------------------------------------------\n");
    $timeformat(-9,0," ns");
    $write("stop time:    %t\n",$stime);
    $write("stop condition: TestBench watchdog\n");
    $write("clk:               %d MHz\n", SYSTEM_CLOCK);
    $write("----------------------------------------------------------------\n");
    $stop(2);
end : stop_WatchDog

//------------------------------------------------------------------------------
always_ff @(posedge clk) begin
    if(rst) begin
        sw <= '0;
    end
    else begin
        sw <= sw + 1'b1;
    end
end

//==============================================================================
//    Instances
//==============================================================================

//------------------------------------------------------------------------------
//    slon5_m
//------------------------------------------------------------------------------

slon5_test slon5
(
    .ref_clk ( clk     ),
    
    .sw      ( sw      ),
             
    .dout    ( dout    ),
    .dnum    ( dnum    )
);

//==============================================================================
//    test & debug
//==============================================================================

//------------------------------------------------------------------------------
initial begin
    $write("----------------------------------------------------------------\n");
    $write("Verify const and parameters\n");
    $write("----------------------------------------------------------------\n");
    $write("\n");
    if(checkKTable(KTable, RefKTable)) begin
        $write("KTable: verify OK!\n");
    end
    else begin
        $error("KTable: verify FAIL!\n");
    end
    $write("\n");
    $write("----------------------------------------------------------------\n");
    $write("end of verification\n");
    $write("----------------------------------------------------------------\n");

    printKTable(KTable);
    printSTable();
    
    $write("WORD_WIDTH:  %2d\n", $clog2(WORD_WIDTH));
    $write("STAGE_WIDTH: %2d\n", $clog2(STAGE_NUM));
end

endmodule : slon5_tb

